module tb_top
(
);

reg [31:0]instruction;
wire [63:0]ReadData1, ReadData2;
  
top t1
(
);

